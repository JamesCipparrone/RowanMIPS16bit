module Register16Bit_tb ();

endmodule
